<<<<<<< HEAD
localparam INDEX_SIZE = 64;
=======
localparam [63:0] INDEX[0:7] = '{ 0, 1, 2, 3, 4, 5, 6, 7 };
>>>>>>> ef81c50a49672289e662a1a1b043a3697a83b61a
