localparam [63:0] INDEX[0:7] = '{ 0, 1, 2, 3, 4, 5, 6, 7 };
