localparam INDEX_SIZE = 64;
